// base_hps.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module base_hps (
		input  wire        clk_clk,                                //                             clk.clk
		input  wire        hps_0_can0_rxd,                         //                      hps_0_can0.rxd
		output wire        hps_0_can0_txd,                         //                                .txd
		output wire [14:0] hps_0_ddr_mem_a,                        //                       hps_0_ddr.mem_a
		output wire [2:0]  hps_0_ddr_mem_ba,                       //                                .mem_ba
		output wire        hps_0_ddr_mem_ck,                       //                                .mem_ck
		output wire        hps_0_ddr_mem_ck_n,                     //                                .mem_ck_n
		output wire        hps_0_ddr_mem_cke,                      //                                .mem_cke
		output wire        hps_0_ddr_mem_cs_n,                     //                                .mem_cs_n
		output wire        hps_0_ddr_mem_ras_n,                    //                                .mem_ras_n
		output wire        hps_0_ddr_mem_cas_n,                    //                                .mem_cas_n
		output wire        hps_0_ddr_mem_we_n,                     //                                .mem_we_n
		output wire        hps_0_ddr_mem_reset_n,                  //                                .mem_reset_n
		inout  wire [31:0] hps_0_ddr_mem_dq,                       //                                .mem_dq
		inout  wire [3:0]  hps_0_ddr_mem_dqs,                      //                                .mem_dqs
		inout  wire [3:0]  hps_0_ddr_mem_dqs_n,                    //                                .mem_dqs_n
		output wire        hps_0_ddr_mem_odt,                      //                                .mem_odt
		output wire [3:0]  hps_0_ddr_mem_dm,                       //                                .mem_dm
		input  wire        hps_0_ddr_oct_rzqin,                    //                                .oct_rzqin
		input  wire [31:0] hps_0_h2f_gp_gp_in,                     //                    hps_0_h2f_gp.gp_in
		output wire [31:0] hps_0_h2f_gp_gp_out,                    //                                .gp_out
		output wire        hps_0_i2c1_out_data,                    //                      hps_0_i2c1.out_data
		input  wire        hps_0_i2c1_sda,                         //                                .sda
		output wire        hps_0_i2c1_clk_clk,                     //                  hps_0_i2c1_clk.clk
		input  wire        hps_0_i2c1_scl_in_clk,                  //               hps_0_i2c1_scl_in.clk
		output wire        hps_0_i2c3_out_data,                    //                      hps_0_i2c3.out_data
		input  wire        hps_0_i2c3_sda,                         //                                .sda
		output wire        hps_0_i2c3_clk_clk,                     //                  hps_0_i2c3_clk.clk
		input  wire        hps_0_i2c3_scl_in_clk,                  //               hps_0_i2c3_scl_in.clk
		output wire        hps_0_io_hps_io_emac1_inst_TX_CLK,      //                        hps_0_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_io_hps_io_emac1_inst_TXD0,        //                                .hps_io_emac1_inst_TXD0
		output wire        hps_0_io_hps_io_emac1_inst_TXD1,        //                                .hps_io_emac1_inst_TXD1
		output wire        hps_0_io_hps_io_emac1_inst_TXD2,        //                                .hps_io_emac1_inst_TXD2
		output wire        hps_0_io_hps_io_emac1_inst_TXD3,        //                                .hps_io_emac1_inst_TXD3
		input  wire        hps_0_io_hps_io_emac1_inst_RXD0,        //                                .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_io_hps_io_emac1_inst_MDIO,        //                                .hps_io_emac1_inst_MDIO
		output wire        hps_0_io_hps_io_emac1_inst_MDC,         //                                .hps_io_emac1_inst_MDC
		input  wire        hps_0_io_hps_io_emac1_inst_RX_CTL,      //                                .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_io_hps_io_emac1_inst_TX_CTL,      //                                .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_io_hps_io_emac1_inst_RX_CLK,      //                                .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_io_hps_io_emac1_inst_RXD1,        //                                .hps_io_emac1_inst_RXD1
		input  wire        hps_0_io_hps_io_emac1_inst_RXD2,        //                                .hps_io_emac1_inst_RXD2
		input  wire        hps_0_io_hps_io_emac1_inst_RXD3,        //                                .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_io_hps_io_sdio_inst_CMD,          //                                .hps_io_sdio_inst_CMD
		inout  wire        hps_0_io_hps_io_sdio_inst_D0,           //                                .hps_io_sdio_inst_D0
		inout  wire        hps_0_io_hps_io_sdio_inst_D1,           //                                .hps_io_sdio_inst_D1
		output wire        hps_0_io_hps_io_sdio_inst_CLK,          //                                .hps_io_sdio_inst_CLK
		inout  wire        hps_0_io_hps_io_sdio_inst_D2,           //                                .hps_io_sdio_inst_D2
		inout  wire        hps_0_io_hps_io_sdio_inst_D3,           //                                .hps_io_sdio_inst_D3
		inout  wire        hps_0_io_hps_io_usb1_inst_D0,           //                                .hps_io_usb1_inst_D0
		inout  wire        hps_0_io_hps_io_usb1_inst_D1,           //                                .hps_io_usb1_inst_D1
		inout  wire        hps_0_io_hps_io_usb1_inst_D2,           //                                .hps_io_usb1_inst_D2
		inout  wire        hps_0_io_hps_io_usb1_inst_D3,           //                                .hps_io_usb1_inst_D3
		inout  wire        hps_0_io_hps_io_usb1_inst_D4,           //                                .hps_io_usb1_inst_D4
		inout  wire        hps_0_io_hps_io_usb1_inst_D5,           //                                .hps_io_usb1_inst_D5
		inout  wire        hps_0_io_hps_io_usb1_inst_D6,           //                                .hps_io_usb1_inst_D6
		inout  wire        hps_0_io_hps_io_usb1_inst_D7,           //                                .hps_io_usb1_inst_D7
		input  wire        hps_0_io_hps_io_usb1_inst_CLK,          //                                .hps_io_usb1_inst_CLK
		output wire        hps_0_io_hps_io_usb1_inst_STP,          //                                .hps_io_usb1_inst_STP
		input  wire        hps_0_io_hps_io_usb1_inst_DIR,          //                                .hps_io_usb1_inst_DIR
		input  wire        hps_0_io_hps_io_usb1_inst_NXT,          //                                .hps_io_usb1_inst_NXT
		input  wire        hps_0_io_hps_io_uart0_inst_RX,          //                                .hps_io_uart0_inst_RX
		output wire        hps_0_io_hps_io_uart0_inst_TX,          //                                .hps_io_uart0_inst_TX
		inout  wire        hps_0_io_hps_io_i2c0_inst_SDA,          //                                .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_io_hps_io_i2c0_inst_SCL,          //                                .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_io_hps_io_gpio_inst_GPIO53,       //                                .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_io_hps_io_gpio_inst_GPIO54,       //                                .hps_io_gpio_inst_GPIO54
		output wire        hps_0_spim0_txd,                        //                     hps_0_spim0.txd
		input  wire        hps_0_spim0_rxd,                        //                                .rxd
		input  wire        hps_0_spim0_ss_in_n,                    //                                .ss_in_n
		output wire        hps_0_spim0_ssi_oe_n,                   //                                .ssi_oe_n
		output wire        hps_0_spim0_ss_0_n,                     //                                .ss_0_n
		output wire        hps_0_spim0_ss_1_n,                     //                                .ss_1_n
		output wire        hps_0_spim0_ss_2_n,                     //                                .ss_2_n
		output wire        hps_0_spim0_ss_3_n,                     //                                .ss_3_n
		output wire        hps_0_spim0_sclk_out_clk,               //            hps_0_spim0_sclk_out.clk
		output wire        hps_0_spim1_txd,                        //                     hps_0_spim1.txd
		input  wire        hps_0_spim1_rxd,                        //                                .rxd
		input  wire        hps_0_spim1_ss_in_n,                    //                                .ss_in_n
		output wire        hps_0_spim1_ssi_oe_n,                   //                                .ssi_oe_n
		output wire        hps_0_spim1_ss_0_n,                     //                                .ss_0_n
		output wire        hps_0_spim1_ss_1_n,                     //                                .ss_1_n
		output wire        hps_0_spim1_ss_2_n,                     //                                .ss_2_n
		output wire        hps_0_spim1_ss_3_n,                     //                                .ss_3_n
		output wire        hps_0_spim1_sclk_out_clk,               //            hps_0_spim1_sclk_out.clk
		input  wire        hps_0_uart1_cts,                        //                     hps_0_uart1.cts
		input  wire        hps_0_uart1_dsr,                        //                                .dsr
		input  wire        hps_0_uart1_dcd,                        //                                .dcd
		input  wire        hps_0_uart1_ri,                         //                                .ri
		output wire        hps_0_uart1_dtr,                        //                                .dtr
		output wire        hps_0_uart1_rts,                        //                                .rts
		output wire        hps_0_uart1_out1_n,                     //                                .out1_n
		output wire        hps_0_uart1_out2_n,                     //                                .out2_n
		input  wire        hps_0_uart1_rxd,                        //                                .rxd
		output wire        hps_0_uart1_txd,                        //                                .txd
		output wire [7:0]  led_pio_external_connection_export,     //     led_pio_external_connection.export
		output wire [8:0]  motor_left_external_connection_export,  //  motor_left_external_connection.export
		output wire [8:0]  motor_right_external_connection_export, // motor_right_external_connection.export
		input  wire [1:0]  pb_pio_external_connection_export,      //      pb_pio_external_connection.export
		output wire        pll_adc_clk_locked_export,              //              pll_adc_clk_locked.export
		output wire        pll_adc_clk_outclk1_clk,                //             pll_adc_clk_outclk1.clk
		input  wire [3:0]  sw_pio_external_connection_export       //      sw_pio_external_connection.export
	);

	wire         hps_0_h2f_cold_reset_reset;                     // hps_0:h2f_cold_rst_n -> [pll_adc_clk:rst, rst_controller:reset_in0]
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                  // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                  // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                 // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                  // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                    // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                 // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                 // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                 // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                 // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                  // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                   // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                 // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                 // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                 // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                 // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                 // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                  // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                   // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                 // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata; // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;  // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_0_led_pio_s1_chipselect;        // mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_0_led_pio_s1_readdata;          // led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_led_pio_s1_address;           // mm_interconnect_0:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_0_led_pio_s1_write;             // mm_interconnect_0:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_0_led_pio_s1_writedata;         // mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	wire  [31:0] mm_interconnect_0_pb_pio_s1_readdata;           // pb_pio:readdata -> mm_interconnect_0:pb_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_pb_pio_s1_address;            // mm_interconnect_0:pb_pio_s1_address -> pb_pio:address
	wire  [31:0] mm_interconnect_0_sw_pio_s1_readdata;           // sw_pio:readdata -> mm_interconnect_0:sw_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_pio_s1_address;            // mm_interconnect_0:sw_pio_s1_address -> sw_pio:address
	wire         mm_interconnect_0_motor_left_s1_chipselect;     // mm_interconnect_0:motor_left_s1_chipselect -> motor_left:chipselect
	wire  [31:0] mm_interconnect_0_motor_left_s1_readdata;       // motor_left:readdata -> mm_interconnect_0:motor_left_s1_readdata
	wire   [1:0] mm_interconnect_0_motor_left_s1_address;        // mm_interconnect_0:motor_left_s1_address -> motor_left:address
	wire         mm_interconnect_0_motor_left_s1_write;          // mm_interconnect_0:motor_left_s1_write -> motor_left:write_n
	wire  [31:0] mm_interconnect_0_motor_left_s1_writedata;      // mm_interconnect_0:motor_left_s1_writedata -> motor_left:writedata
	wire         mm_interconnect_0_motor_right_s1_chipselect;    // mm_interconnect_0:motor_right_s1_chipselect -> motor_right:chipselect
	wire  [31:0] mm_interconnect_0_motor_right_s1_readdata;      // motor_right:readdata -> mm_interconnect_0:motor_right_s1_readdata
	wire   [1:0] mm_interconnect_0_motor_right_s1_address;       // mm_interconnect_0:motor_right_s1_address -> motor_right:address
	wire         mm_interconnect_0_motor_right_s1_write;         // mm_interconnect_0:motor_right_s1_write -> motor_right:write_n
	wire  [31:0] mm_interconnect_0_motor_right_s1_writedata;     // mm_interconnect_0:motor_right_s1_writedata -> motor_right:writedata
	wire         rst_controller_reset_out_reset;                 // rst_controller:reset_out -> [led_pio:reset_n, mm_interconnect_0:sysid_reset_reset_bridge_in_reset_reset, pb_pio:reset_n, sw_pio:reset_n, sysid:reset_n]
	wire         hps_0_h2f_reset_reset;                          // hps_0:h2f_rst_n -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;             // rst_controller_001:reset_out -> [mm_interconnect_0:motor_left_reset_reset_bridge_in_reset_reset, motor_left:reset_n, motor_right:reset_n]

	base_hps_hps_0 #(
		.F2S_Width (1),
		.S2F_Width (1)
	) hps_0 (
		.h2f_cold_rst_n           (hps_0_h2f_cold_reset_reset),        //           h2f_cold_reset.reset_n
		.h2f_pending_rst_req_n    (),                                  // h2f_warm_reset_handshake.h2f_pending_rst_req_n
		.f2h_pending_rst_ack_n    (),                                  //                         .f2h_pending_rst_ack_n
		.h2f_gp_in                (hps_0_h2f_gp_gp_in),                //                   h2f_gp.gp_in
		.h2f_gp_out               (hps_0_h2f_gp_gp_out),               //                         .gp_out
		.spim0_txd                (hps_0_spim0_txd),                   //                    spim0.txd
		.spim0_rxd                (hps_0_spim0_rxd),                   //                         .rxd
		.spim0_ss_in_n            (hps_0_spim0_ss_in_n),               //                         .ss_in_n
		.spim0_ssi_oe_n           (hps_0_spim0_ssi_oe_n),              //                         .ssi_oe_n
		.spim0_ss_0_n             (hps_0_spim0_ss_0_n),                //                         .ss_0_n
		.spim0_ss_1_n             (hps_0_spim0_ss_1_n),                //                         .ss_1_n
		.spim0_ss_2_n             (hps_0_spim0_ss_2_n),                //                         .ss_2_n
		.spim0_ss_3_n             (hps_0_spim0_ss_3_n),                //                         .ss_3_n
		.spim0_sclk_out           (hps_0_spim0_sclk_out_clk),          //           spim0_sclk_out.clk
		.spim1_txd                (hps_0_spim1_txd),                   //                    spim1.txd
		.spim1_rxd                (hps_0_spim1_rxd),                   //                         .rxd
		.spim1_ss_in_n            (hps_0_spim1_ss_in_n),               //                         .ss_in_n
		.spim1_ssi_oe_n           (hps_0_spim1_ssi_oe_n),              //                         .ssi_oe_n
		.spim1_ss_0_n             (hps_0_spim1_ss_0_n),                //                         .ss_0_n
		.spim1_ss_1_n             (hps_0_spim1_ss_1_n),                //                         .ss_1_n
		.spim1_ss_2_n             (hps_0_spim1_ss_2_n),                //                         .ss_2_n
		.spim1_ss_3_n             (hps_0_spim1_ss_3_n),                //                         .ss_3_n
		.spim1_sclk_out           (hps_0_spim1_sclk_out_clk),          //           spim1_sclk_out.clk
		.uart1_cts                (hps_0_uart1_cts),                   //                    uart1.cts
		.uart1_dsr                (hps_0_uart1_dsr),                   //                         .dsr
		.uart1_dcd                (hps_0_uart1_dcd),                   //                         .dcd
		.uart1_ri                 (hps_0_uart1_ri),                    //                         .ri
		.uart1_dtr                (hps_0_uart1_dtr),                   //                         .dtr
		.uart1_rts                (hps_0_uart1_rts),                   //                         .rts
		.uart1_out1_n             (hps_0_uart1_out1_n),                //                         .out1_n
		.uart1_out2_n             (hps_0_uart1_out2_n),                //                         .out2_n
		.uart1_rxd                (hps_0_uart1_rxd),                   //                         .rxd
		.uart1_txd                (hps_0_uart1_txd),                   //                         .txd
		.i2c1_scl                 (hps_0_i2c1_scl_in_clk),             //              i2c1_scl_in.clk
		.i2c1_out_clk             (hps_0_i2c1_clk_clk),                //                 i2c1_clk.clk
		.i2c1_out_data            (hps_0_i2c1_out_data),               //                     i2c1.out_data
		.i2c1_sda                 (hps_0_i2c1_sda),                    //                         .sda
		.i2c_emac1_scl            (hps_0_i2c3_scl_in_clk),             //              i2c3_scl_in.clk
		.i2c_emac1_out_clk        (hps_0_i2c3_clk_clk),                //                 i2c3_clk.clk
		.i2c_emac1_out_data       (hps_0_i2c3_out_data),               //                     i2c3.out_data
		.i2c_emac1_sda            (hps_0_i2c3_sda),                    //                         .sda
		.can0_rxd                 (hps_0_can0_rxd),                    //                     can0.rxd
		.can0_txd                 (hps_0_can0_txd),                    //                         .txd
		.mem_a                    (hps_0_ddr_mem_a),                   //                   memory.mem_a
		.mem_ba                   (hps_0_ddr_mem_ba),                  //                         .mem_ba
		.mem_ck                   (hps_0_ddr_mem_ck),                  //                         .mem_ck
		.mem_ck_n                 (hps_0_ddr_mem_ck_n),                //                         .mem_ck_n
		.mem_cke                  (hps_0_ddr_mem_cke),                 //                         .mem_cke
		.mem_cs_n                 (hps_0_ddr_mem_cs_n),                //                         .mem_cs_n
		.mem_ras_n                (hps_0_ddr_mem_ras_n),               //                         .mem_ras_n
		.mem_cas_n                (hps_0_ddr_mem_cas_n),               //                         .mem_cas_n
		.mem_we_n                 (hps_0_ddr_mem_we_n),                //                         .mem_we_n
		.mem_reset_n              (hps_0_ddr_mem_reset_n),             //                         .mem_reset_n
		.mem_dq                   (hps_0_ddr_mem_dq),                  //                         .mem_dq
		.mem_dqs                  (hps_0_ddr_mem_dqs),                 //                         .mem_dqs
		.mem_dqs_n                (hps_0_ddr_mem_dqs_n),               //                         .mem_dqs_n
		.mem_odt                  (hps_0_ddr_mem_odt),                 //                         .mem_odt
		.mem_dm                   (hps_0_ddr_mem_dm),                  //                         .mem_dm
		.oct_rzqin                (hps_0_ddr_oct_rzqin),               //                         .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_io_hps_io_emac1_inst_TX_CLK), //                   hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_io_hps_io_emac1_inst_TXD0),   //                         .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_io_hps_io_emac1_inst_TXD1),   //                         .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_io_hps_io_emac1_inst_TXD2),   //                         .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_io_hps_io_emac1_inst_TXD3),   //                         .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_io_hps_io_emac1_inst_RXD0),   //                         .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_io_hps_io_emac1_inst_MDIO),   //                         .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_io_hps_io_emac1_inst_MDC),    //                         .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_io_hps_io_emac1_inst_RX_CTL), //                         .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_io_hps_io_emac1_inst_TX_CTL), //                         .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_io_hps_io_emac1_inst_RX_CLK), //                         .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_io_hps_io_emac1_inst_RXD1),   //                         .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_io_hps_io_emac1_inst_RXD2),   //                         .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_io_hps_io_emac1_inst_RXD3),   //                         .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_0_io_hps_io_sdio_inst_CMD),     //                         .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_io_hps_io_sdio_inst_D0),      //                         .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_io_hps_io_sdio_inst_D1),      //                         .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_io_hps_io_sdio_inst_CLK),     //                         .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_io_hps_io_sdio_inst_D2),      //                         .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_io_hps_io_sdio_inst_D3),      //                         .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_io_hps_io_usb1_inst_D0),      //                         .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_io_hps_io_usb1_inst_D1),      //                         .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_io_hps_io_usb1_inst_D2),      //                         .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_io_hps_io_usb1_inst_D3),      //                         .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_io_hps_io_usb1_inst_D4),      //                         .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_io_hps_io_usb1_inst_D5),      //                         .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_io_hps_io_usb1_inst_D6),      //                         .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_io_hps_io_usb1_inst_D7),      //                         .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_io_hps_io_usb1_inst_CLK),     //                         .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_io_hps_io_usb1_inst_STP),     //                         .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_io_hps_io_usb1_inst_DIR),     //                         .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_io_hps_io_usb1_inst_NXT),     //                         .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (hps_0_io_hps_io_uart0_inst_RX),     //                         .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_io_hps_io_uart0_inst_TX),     //                         .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_io_hps_io_i2c0_inst_SDA),     //                         .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_io_hps_io_i2c0_inst_SCL),     //                         .hps_io_i2c0_inst_SCL
		.hps_io_gpio_inst_GPIO53  (hps_0_io_hps_io_gpio_inst_GPIO53),  //                         .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_io_hps_io_gpio_inst_GPIO54),  //                         .hps_io_gpio_inst_GPIO54
		.h2f_rst_n                (hps_0_h2f_reset_reset),             //                h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                           //            h2f_axi_clock.clk
		.h2f_AWID                 (),                                  //           h2f_axi_master.awid
		.h2f_AWADDR               (),                                  //                         .awaddr
		.h2f_AWLEN                (),                                  //                         .awlen
		.h2f_AWSIZE               (),                                  //                         .awsize
		.h2f_AWBURST              (),                                  //                         .awburst
		.h2f_AWLOCK               (),                                  //                         .awlock
		.h2f_AWCACHE              (),                                  //                         .awcache
		.h2f_AWPROT               (),                                  //                         .awprot
		.h2f_AWVALID              (),                                  //                         .awvalid
		.h2f_AWREADY              (),                                  //                         .awready
		.h2f_WID                  (),                                  //                         .wid
		.h2f_WDATA                (),                                  //                         .wdata
		.h2f_WSTRB                (),                                  //                         .wstrb
		.h2f_WLAST                (),                                  //                         .wlast
		.h2f_WVALID               (),                                  //                         .wvalid
		.h2f_WREADY               (),                                  //                         .wready
		.h2f_BID                  (),                                  //                         .bid
		.h2f_BRESP                (),                                  //                         .bresp
		.h2f_BVALID               (),                                  //                         .bvalid
		.h2f_BREADY               (),                                  //                         .bready
		.h2f_ARID                 (),                                  //                         .arid
		.h2f_ARADDR               (),                                  //                         .araddr
		.h2f_ARLEN                (),                                  //                         .arlen
		.h2f_ARSIZE               (),                                  //                         .arsize
		.h2f_ARBURST              (),                                  //                         .arburst
		.h2f_ARLOCK               (),                                  //                         .arlock
		.h2f_ARCACHE              (),                                  //                         .arcache
		.h2f_ARPROT               (),                                  //                         .arprot
		.h2f_ARVALID              (),                                  //                         .arvalid
		.h2f_ARREADY              (),                                  //                         .arready
		.h2f_RID                  (),                                  //                         .rid
		.h2f_RDATA                (),                                  //                         .rdata
		.h2f_RRESP                (),                                  //                         .rresp
		.h2f_RLAST                (),                                  //                         .rlast
		.h2f_RVALID               (),                                  //                         .rvalid
		.h2f_RREADY               (),                                  //                         .rready
		.f2h_axi_clk              (clk_clk),                           //            f2h_axi_clock.clk
		.f2h_AWID                 (),                                  //            f2h_axi_slave.awid
		.f2h_AWADDR               (),                                  //                         .awaddr
		.f2h_AWLEN                (),                                  //                         .awlen
		.f2h_AWSIZE               (),                                  //                         .awsize
		.f2h_AWBURST              (),                                  //                         .awburst
		.f2h_AWLOCK               (),                                  //                         .awlock
		.f2h_AWCACHE              (),                                  //                         .awcache
		.f2h_AWPROT               (),                                  //                         .awprot
		.f2h_AWVALID              (),                                  //                         .awvalid
		.f2h_AWREADY              (),                                  //                         .awready
		.f2h_AWUSER               (),                                  //                         .awuser
		.f2h_WID                  (),                                  //                         .wid
		.f2h_WDATA                (),                                  //                         .wdata
		.f2h_WSTRB                (),                                  //                         .wstrb
		.f2h_WLAST                (),                                  //                         .wlast
		.f2h_WVALID               (),                                  //                         .wvalid
		.f2h_WREADY               (),                                  //                         .wready
		.f2h_BID                  (),                                  //                         .bid
		.f2h_BRESP                (),                                  //                         .bresp
		.f2h_BVALID               (),                                  //                         .bvalid
		.f2h_BREADY               (),                                  //                         .bready
		.f2h_ARID                 (),                                  //                         .arid
		.f2h_ARADDR               (),                                  //                         .araddr
		.f2h_ARLEN                (),                                  //                         .arlen
		.f2h_ARSIZE               (),                                  //                         .arsize
		.f2h_ARBURST              (),                                  //                         .arburst
		.f2h_ARLOCK               (),                                  //                         .arlock
		.f2h_ARCACHE              (),                                  //                         .arcache
		.f2h_ARPROT               (),                                  //                         .arprot
		.f2h_ARVALID              (),                                  //                         .arvalid
		.f2h_ARREADY              (),                                  //                         .arready
		.f2h_ARUSER               (),                                  //                         .aruser
		.f2h_RID                  (),                                  //                         .rid
		.f2h_RDATA                (),                                  //                         .rdata
		.f2h_RRESP                (),                                  //                         .rresp
		.f2h_RLAST                (),                                  //                         .rlast
		.f2h_RVALID               (),                                  //                         .rvalid
		.f2h_RREADY               (),                                  //                         .rready
		.h2f_lw_axi_clk           (clk_clk),                           //         h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),      //        h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),    //                         .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),     //                         .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),    //                         .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),   //                         .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),    //                         .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),   //                         .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),    //                         .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),   //                         .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),   //                         .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),       //                         .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),     //                         .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),     //                         .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),     //                         .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),    //                         .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),    //                         .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),       //                         .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),     //                         .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),    //                         .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),    //                         .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),      //                         .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),    //                         .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),     //                         .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),    //                         .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),   //                         .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),    //                         .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),   //                         .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),    //                         .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),   //                         .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),   //                         .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),       //                         .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),     //                         .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),     //                         .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),     //                         .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),    //                         .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)     //                         .rready
	);

	base_hps_led_pio led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)       // external_connection.export
	);

	base_hps_motor_left motor_left (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_motor_left_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_motor_left_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_motor_left_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_motor_left_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_motor_left_s1_readdata),   //                    .readdata
		.out_port   (motor_left_external_connection_export)       // external_connection.export
	);

	base_hps_motor_left motor_right (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_motor_right_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_motor_right_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_motor_right_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_motor_right_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_motor_right_s1_readdata),   //                    .readdata
		.out_port   (motor_right_external_connection_export)       // external_connection.export
	);

	base_hps_pb_pio pb_pio (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_pb_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pb_pio_s1_readdata), //                    .readdata
		.in_port  (pb_pio_external_connection_export)     // external_connection.export
	);

	base_hps_pll_adc_clk pll_adc_clk (
		.refclk   (clk_clk),                     //  refclk.clk
		.rst      (~hps_0_h2f_cold_reset_reset), //   reset.reset
		.outclk_0 (),                            // outclk0.clk
		.outclk_1 (pll_adc_clk_outclk1_clk),     // outclk1.clk
		.locked   (pll_adc_clk_locked_export)    //  locked.export
	);

	base_hps_sw_pio sw_pio (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_sw_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_pio_s1_readdata), //                    .readdata
		.in_port  (sw_pio_external_connection_export)     // external_connection.export
	);

	base_hps_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	base_hps_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                 (hps_0_h2f_lw_axi_master_awid),                   //                hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr               (hps_0_h2f_lw_axi_master_awaddr),                 //                                       .awaddr
		.hps_0_h2f_lw_axi_master_awlen                (hps_0_h2f_lw_axi_master_awlen),                  //                                       .awlen
		.hps_0_h2f_lw_axi_master_awsize               (hps_0_h2f_lw_axi_master_awsize),                 //                                       .awsize
		.hps_0_h2f_lw_axi_master_awburst              (hps_0_h2f_lw_axi_master_awburst),                //                                       .awburst
		.hps_0_h2f_lw_axi_master_awlock               (hps_0_h2f_lw_axi_master_awlock),                 //                                       .awlock
		.hps_0_h2f_lw_axi_master_awcache              (hps_0_h2f_lw_axi_master_awcache),                //                                       .awcache
		.hps_0_h2f_lw_axi_master_awprot               (hps_0_h2f_lw_axi_master_awprot),                 //                                       .awprot
		.hps_0_h2f_lw_axi_master_awvalid              (hps_0_h2f_lw_axi_master_awvalid),                //                                       .awvalid
		.hps_0_h2f_lw_axi_master_awready              (hps_0_h2f_lw_axi_master_awready),                //                                       .awready
		.hps_0_h2f_lw_axi_master_wid                  (hps_0_h2f_lw_axi_master_wid),                    //                                       .wid
		.hps_0_h2f_lw_axi_master_wdata                (hps_0_h2f_lw_axi_master_wdata),                  //                                       .wdata
		.hps_0_h2f_lw_axi_master_wstrb                (hps_0_h2f_lw_axi_master_wstrb),                  //                                       .wstrb
		.hps_0_h2f_lw_axi_master_wlast                (hps_0_h2f_lw_axi_master_wlast),                  //                                       .wlast
		.hps_0_h2f_lw_axi_master_wvalid               (hps_0_h2f_lw_axi_master_wvalid),                 //                                       .wvalid
		.hps_0_h2f_lw_axi_master_wready               (hps_0_h2f_lw_axi_master_wready),                 //                                       .wready
		.hps_0_h2f_lw_axi_master_bid                  (hps_0_h2f_lw_axi_master_bid),                    //                                       .bid
		.hps_0_h2f_lw_axi_master_bresp                (hps_0_h2f_lw_axi_master_bresp),                  //                                       .bresp
		.hps_0_h2f_lw_axi_master_bvalid               (hps_0_h2f_lw_axi_master_bvalid),                 //                                       .bvalid
		.hps_0_h2f_lw_axi_master_bready               (hps_0_h2f_lw_axi_master_bready),                 //                                       .bready
		.hps_0_h2f_lw_axi_master_arid                 (hps_0_h2f_lw_axi_master_arid),                   //                                       .arid
		.hps_0_h2f_lw_axi_master_araddr               (hps_0_h2f_lw_axi_master_araddr),                 //                                       .araddr
		.hps_0_h2f_lw_axi_master_arlen                (hps_0_h2f_lw_axi_master_arlen),                  //                                       .arlen
		.hps_0_h2f_lw_axi_master_arsize               (hps_0_h2f_lw_axi_master_arsize),                 //                                       .arsize
		.hps_0_h2f_lw_axi_master_arburst              (hps_0_h2f_lw_axi_master_arburst),                //                                       .arburst
		.hps_0_h2f_lw_axi_master_arlock               (hps_0_h2f_lw_axi_master_arlock),                 //                                       .arlock
		.hps_0_h2f_lw_axi_master_arcache              (hps_0_h2f_lw_axi_master_arcache),                //                                       .arcache
		.hps_0_h2f_lw_axi_master_arprot               (hps_0_h2f_lw_axi_master_arprot),                 //                                       .arprot
		.hps_0_h2f_lw_axi_master_arvalid              (hps_0_h2f_lw_axi_master_arvalid),                //                                       .arvalid
		.hps_0_h2f_lw_axi_master_arready              (hps_0_h2f_lw_axi_master_arready),                //                                       .arready
		.hps_0_h2f_lw_axi_master_rid                  (hps_0_h2f_lw_axi_master_rid),                    //                                       .rid
		.hps_0_h2f_lw_axi_master_rdata                (hps_0_h2f_lw_axi_master_rdata),                  //                                       .rdata
		.hps_0_h2f_lw_axi_master_rresp                (hps_0_h2f_lw_axi_master_rresp),                  //                                       .rresp
		.hps_0_h2f_lw_axi_master_rlast                (hps_0_h2f_lw_axi_master_rlast),                  //                                       .rlast
		.hps_0_h2f_lw_axi_master_rvalid               (hps_0_h2f_lw_axi_master_rvalid),                 //                                       .rvalid
		.hps_0_h2f_lw_axi_master_rready               (hps_0_h2f_lw_axi_master_rready),                 //                                       .rready
		.clk_0_clk_clk                                (clk_clk),                                        //                              clk_0_clk.clk
		.motor_left_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),             // motor_left_reset_reset_bridge_in_reset.reset
		.sysid_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                 //      sysid_reset_reset_bridge_in_reset.reset
		.led_pio_s1_address                           (mm_interconnect_0_led_pio_s1_address),           //                             led_pio_s1.address
		.led_pio_s1_write                             (mm_interconnect_0_led_pio_s1_write),             //                                       .write
		.led_pio_s1_readdata                          (mm_interconnect_0_led_pio_s1_readdata),          //                                       .readdata
		.led_pio_s1_writedata                         (mm_interconnect_0_led_pio_s1_writedata),         //                                       .writedata
		.led_pio_s1_chipselect                        (mm_interconnect_0_led_pio_s1_chipselect),        //                                       .chipselect
		.motor_left_s1_address                        (mm_interconnect_0_motor_left_s1_address),        //                          motor_left_s1.address
		.motor_left_s1_write                          (mm_interconnect_0_motor_left_s1_write),          //                                       .write
		.motor_left_s1_readdata                       (mm_interconnect_0_motor_left_s1_readdata),       //                                       .readdata
		.motor_left_s1_writedata                      (mm_interconnect_0_motor_left_s1_writedata),      //                                       .writedata
		.motor_left_s1_chipselect                     (mm_interconnect_0_motor_left_s1_chipselect),     //                                       .chipselect
		.motor_right_s1_address                       (mm_interconnect_0_motor_right_s1_address),       //                         motor_right_s1.address
		.motor_right_s1_write                         (mm_interconnect_0_motor_right_s1_write),         //                                       .write
		.motor_right_s1_readdata                      (mm_interconnect_0_motor_right_s1_readdata),      //                                       .readdata
		.motor_right_s1_writedata                     (mm_interconnect_0_motor_right_s1_writedata),     //                                       .writedata
		.motor_right_s1_chipselect                    (mm_interconnect_0_motor_right_s1_chipselect),    //                                       .chipselect
		.pb_pio_s1_address                            (mm_interconnect_0_pb_pio_s1_address),            //                              pb_pio_s1.address
		.pb_pio_s1_readdata                           (mm_interconnect_0_pb_pio_s1_readdata),           //                                       .readdata
		.sw_pio_s1_address                            (mm_interconnect_0_sw_pio_s1_address),            //                              sw_pio_s1.address
		.sw_pio_s1_readdata                           (mm_interconnect_0_sw_pio_s1_readdata),           //                                       .readdata
		.sysid_control_slave_address                  (mm_interconnect_0_sysid_control_slave_address),  //                    sysid_control_slave.address
		.sysid_control_slave_readdata                 (mm_interconnect_0_sysid_control_slave_readdata)  //                                       .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_cold_reset_reset),    // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),         // reset_in1.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
